*charge pump circuit

VDD 1 0 DC 1.20
Vclock1 7 0 DC 0 PULSE(0.00 5.00 1.00N 0.10N 0.10N 1.00N 2.20N)
V14 14 0 DC 1.80V

* Switch Transistors
MN1 7 16 9 0 N1  W= 0.30U L= 0.10U
MN2 7 17 8 0 N1  W= 0.30U L= 0.10U
MN3 7 7 13 0 N1  W= 0.30U L= 0.10U
MN4 7 18 10 0 N1  W= 0.30U L= 0.10U
MN5 14 14 7 0 N1  W= 0.30U L= 0.10U
MN6 14 11 7 0 N1  W= 0.30U L= 0.10U
MN7 14 19 11 0 N1  W= 0.30U L= 0.10U
MN8 0 7 7 0 N1  W= 0.50U L= 0.10U
MP1 8 17 7 1 P1  W= 0.30U L= 0.10U
MP2 9 16 7 1 P1  W= 0.30U L= 0.10U
MP3 10 18 7 1 P1  W= 0.30U L= 0.10U
MP4 11 19 7 1 P1  W= 0.30U L= 0.10U
MP5 1 7 7 1 P1  W= 0.50U L= 0.10U

* charge-transfer capacitors
C1 13 0 10pF
C2 7 0 10pF
C3 7 0 10pF
C4 7 0 10pF
C5 7 0 10pF
C6 7 0 10pF


* n-MOS low leakage
.MODEL N1 NMOS LEVEL=14 VTHO=0.28 U0=0.060 TOXE= 1.2E-9 LINT=0.015U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.570 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  0.9 U0=0.060 UA=3.400e-15
+WINT=0.005U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.010
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p


* p-MOS low leakage
.MODEL P1 PMOS LEVEL=14 VTHO=-0.32 U0=0.027 TOXE= 1.2E-9 LINT=0.015U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.570 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.9 U0=0.027 UA=2.200e-15
+WINT=0.005U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.010
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p


* Transient analysis

.control
tran 0.1N 50.00N
print  V(13) V(7) V(14)
plot  V(13) V(7) V(14)
.endc
.END
